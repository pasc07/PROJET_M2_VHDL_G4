-- mon_sopc.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mon_sopc is
	port (
		avalon_bouton_0_conduit_end_bp_babord       : in  std_logic                    := '0';             -- avalon_bouton_0_conduit_end.bp_babord
		avalon_bouton_0_conduit_end_bp_tribord      : in  std_logic                    := '0';             --                            .bp_tribord
		avalon_bouton_0_conduit_end_bp_stby         : in  std_logic                    := '0';             --                            .bp_stby
		avalon_bouton_0_conduit_end_ledbabord       : out std_logic;                                       --                            .ledbabord
		avalon_bouton_0_conduit_end_ledtribord      : out std_logic;                                       --                            .ledtribord
		avalon_bouton_0_conduit_end_ledstby         : out std_logic;                                       --                            .ledstby
		avalon_bouton_0_conduit_end_out_bip         : out std_logic;                                       --                            .out_bip
		avalon_verin_0_conduit_end_sck_o            : out std_logic;                                       --  avalon_verin_0_conduit_end.sck_o
		avalon_verin_0_conduit_end_pwm_o            : out std_logic;                                       --                            .pwm_o
		avalon_verin_0_conduit_end_sens_o           : out std_logic;                                       --                            .sens_o
		avalon_verin_0_conduit_end_miso_i           : in  std_logic                    := '0';             --                            .miso_i
		avalon_verin_0_conduit_end_cs_n_o           : out std_logic;                                       --                            .cs_n_o
		boutons_external_connection_export          : in  std_logic_vector(1 downto 0) := (others => '0'); -- boutons_external_connection.export
		clk_clk                                     : in  std_logic                    := '0';             --                         clk.clk
		leds_external_connection_export             : out std_logic_vector(7 downto 0);                    --    leds_external_connection.export
		test_anemo_0_conduit_end_beginbursttransfer : in  std_logic                    := '0';             --    test_anemo_0_conduit_end.beginbursttransfer
		test_pwm_0_conduit_end_writeresponsevalid_n : out std_logic                                        --      test_pwm_0_conduit_end.writeresponsevalid_n
	);
end entity mon_sopc;

architecture rtl of mon_sopc is
	component avalon_gestion_bouton is
		port (
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			clk_50M    : in  std_logic                     := 'X';             -- clk
			BP_Babord  : in  std_logic                     := 'X';             -- bp_babord
			BP_Tribord : in  std_logic                     := 'X';             -- bp_tribord
			BP_STBY    : in  std_logic                     := 'X';             -- bp_stby
			ledBabord  : out std_logic;                                        -- ledbabord
			ledTribord : out std_logic;                                        -- ledtribord
			ledSTBY    : out std_logic;                                        -- ledstby
			out_bip    : out std_logic                                         -- out_bip
		);
	end component avalon_gestion_bouton;

	component avalon_verin is
		port (
			write_data_i : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read_data_o  : out std_logic_vector(31 downto 0);                    -- readdata
			address_i    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_i      : in  std_logic                     := 'X';             -- write
			read_i       : in  std_logic                     := 'X';             -- read
			sck_o        : out std_logic;                                        -- sck_o
			pwm_o        : out std_logic;                                        -- pwm_o
			sens_o       : out std_logic;                                        -- sens_o
			miso_i       : in  std_logic                     := 'X';             -- miso_i
			cs_n_o       : out std_logic;                                        -- cs_n_o
			clk_i        : in  std_logic                     := 'X';             -- clk
			arst_i       : in  std_logic                     := 'X'              -- reset
		);
	end component avalon_verin;

	component mon_sopc_boutons is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component mon_sopc_boutons;

	component mon_sopc_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component mon_sopc_jtag_uart_0;

	component mon_sopc_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component mon_sopc_leds;

	component mon_sopc_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component mon_sopc_nios2_gen2_0;

	component mon_sopc_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component mon_sopc_ram;

	component avalon_gestion_anemometre is
		port (
			chipselect         : in  std_logic                     := 'X';             -- chipselect
			write_n            : in  std_logic                     := 'X';             -- write_n
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			clk_50M            : in  std_logic                     := 'X';             -- clk
			in_freq_anemometre : in  std_logic                     := 'X'              -- beginbursttransfer
		);
	end component avalon_gestion_anemometre;

	component avalon_pwm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			out_pwm    : out std_logic                                         -- writeresponsevalid_n
		);
	end component avalon_pwm;

	component mon_sopc_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_bouton_0_avalon_slave_0_address         : out std_logic_vector(1 downto 0);                     -- address
			avalon_bouton_0_avalon_slave_0_write           : out std_logic;                                        -- write
			avalon_bouton_0_avalon_slave_0_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_bouton_0_avalon_slave_0_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_bouton_0_avalon_slave_0_chipselect      : out std_logic;                                        -- chipselect
			avalon_verin_0_avalon_slave_0_address          : out std_logic_vector(2 downto 0);                     -- address
			avalon_verin_0_avalon_slave_0_write            : out std_logic;                                        -- write
			avalon_verin_0_avalon_slave_0_read             : out std_logic;                                        -- read
			avalon_verin_0_avalon_slave_0_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_verin_0_avalon_slave_0_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			boutons_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			boutons_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			leds_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                  : out std_logic;                                        -- write
			leds_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                             : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			ram_s1_address                                 : out std_logic_vector(12 downto 0);                    -- address
			ram_s1_write                                   : out std_logic;                                        -- write
			ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			ram_s1_clken                                   : out std_logic;                                        -- clken
			test_anemo_0_avalon_slave_0_address            : out std_logic_vector(1 downto 0);                     -- address
			test_anemo_0_avalon_slave_0_write              : out std_logic;                                        -- write
			test_anemo_0_avalon_slave_0_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_anemo_0_avalon_slave_0_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			test_anemo_0_avalon_slave_0_chipselect         : out std_logic;                                        -- chipselect
			test_pwm_0_avalon_slave_0_address              : out std_logic_vector(1 downto 0);                     -- address
			test_pwm_0_avalon_slave_0_write                : out std_logic;                                        -- write
			test_pwm_0_avalon_slave_0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_pwm_0_avalon_slave_0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			test_pwm_0_avalon_slave_0_chipselect           : out std_logic                                         -- chipselect
		);
	end component mon_sopc_mm_interconnect_0;

	component mon_sopc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component mon_sopc_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_debug_reset_request_reset                           : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal nios2_gen2_0_data_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                             : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                 : std_logic_vector(16 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                              : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                    : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                   : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                               : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                          : std_logic_vector(16 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                             : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect       : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata         : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest      : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read             : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:test_pwm_0_avalon_slave_0_chipselect -> test_pwm_0:chipselect
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0); -- test_pwm_0:readdata -> mm_interconnect_0:test_pwm_0_avalon_slave_0_readdata
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:test_pwm_0_avalon_slave_0_address -> test_pwm_0:address
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_write                : std_logic;                     -- mm_interconnect_0:test_pwm_0_avalon_slave_0_write -> mm_interconnect_0_test_pwm_0_avalon_slave_0_write:in
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:test_pwm_0_avalon_slave_0_writedata -> test_pwm_0:writedata
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_chipselect         : std_logic;                     -- mm_interconnect_0:test_anemo_0_avalon_slave_0_chipselect -> test_anemo_0:chipselect
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_readdata           : std_logic_vector(31 downto 0); -- test_anemo_0:readdata -> mm_interconnect_0:test_anemo_0_avalon_slave_0_readdata
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:test_anemo_0_avalon_slave_0_address -> test_anemo_0:address
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_write              : std_logic;                     -- mm_interconnect_0:test_anemo_0_avalon_slave_0_write -> mm_interconnect_0_test_anemo_0_avalon_slave_0_write:in
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:test_anemo_0_avalon_slave_0_writedata -> test_anemo_0:writedata
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_chipselect      : std_logic;                     -- mm_interconnect_0:avalon_bouton_0_avalon_slave_0_chipselect -> avalon_bouton_0:chipselect
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- avalon_bouton_0:readdata -> mm_interconnect_0:avalon_bouton_0_avalon_slave_0_readdata
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:avalon_bouton_0_avalon_slave_0_address -> avalon_bouton_0:address
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:avalon_bouton_0_avalon_slave_0_write -> mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write:in
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:avalon_bouton_0_avalon_slave_0_writedata -> avalon_bouton_0:writedata
	signal mm_interconnect_0_avalon_verin_0_avalon_slave_0_readdata         : std_logic_vector(31 downto 0); -- avalon_verin_0:read_data_o -> mm_interconnect_0:avalon_verin_0_avalon_slave_0_readdata
	signal mm_interconnect_0_avalon_verin_0_avalon_slave_0_address          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:avalon_verin_0_avalon_slave_0_address -> avalon_verin_0:address_i
	signal mm_interconnect_0_avalon_verin_0_avalon_slave_0_read             : std_logic;                     -- mm_interconnect_0:avalon_verin_0_avalon_slave_0_read -> avalon_verin_0:read_i
	signal mm_interconnect_0_avalon_verin_0_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:avalon_verin_0_avalon_slave_0_write -> avalon_verin_0:write_i
	signal mm_interconnect_0_avalon_verin_0_avalon_slave_0_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:avalon_verin_0_avalon_slave_0_writedata -> avalon_verin_0:write_data_i
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata          : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest       : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_ram_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	signal mm_interconnect_0_ram_s1_readdata                                : std_logic_vector(31 downto 0); -- ram:readdata -> mm_interconnect_0:ram_s1_readdata
	signal mm_interconnect_0_ram_s1_address                                 : std_logic_vector(12 downto 0); -- mm_interconnect_0:ram_s1_address -> ram:address
	signal mm_interconnect_0_ram_s1_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	signal mm_interconnect_0_ram_s1_write                                   : std_logic;                     -- mm_interconnect_0:ram_s1_write -> ram:write
	signal mm_interconnect_0_ram_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ram_s1_writedata -> ram:writedata
	signal mm_interconnect_0_ram_s1_clken                                   : std_logic;                     -- mm_interconnect_0:ram_s1_clken -> ram:clken
	signal mm_interconnect_0_leds_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                               : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                  : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_boutons_s1_readdata                            : std_logic_vector(31 downto 0); -- boutons:readdata -> mm_interconnect_0:boutons_s1_readdata
	signal mm_interconnect_0_boutons_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:boutons_s1_address -> boutons:address
	signal irq_mapper_receiver0_irq                                         : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                   : std_logic;                     -- rst_controller:reset_out -> [avalon_verin_0:arst_i, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                               : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, ram:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_test_pwm_0_avalon_slave_0_write_ports_inv      : std_logic;                     -- mm_interconnect_0_test_pwm_0_avalon_slave_0_write:inv -> test_pwm_0:write_n
	signal mm_interconnect_0_test_anemo_0_avalon_slave_0_write_ports_inv    : std_logic;                     -- mm_interconnect_0_test_anemo_0_avalon_slave_0_write:inv -> test_anemo_0:write_n
	signal mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write:inv -> avalon_bouton_0:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_reset_out_reset:inv -> [avalon_bouton_0:reset_n, boutons:reset_n, jtag_uart_0:rst_n, leds:reset_n, nios2_gen2_0:reset_n, test_anemo_0:reset_n, test_pwm_0:reset_n]

begin

	avalon_bouton_0 : component avalon_gestion_bouton
		port map (
			chipselect => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_chipselect,      -- avalon_slave_0.chipselect
			write_n    => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write_ports_inv, --               .write_n
			writedata  => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_writedata,       --               .writedata
			readdata   => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_readdata,        --               .readdata
			address    => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_address,         --               .address
			reset_n    => rst_controller_reset_out_reset_ports_inv,                         --          reset.reset_n
			clk_50M    => clk_clk,                                                          --     clock_sink.clk
			BP_Babord  => avalon_bouton_0_conduit_end_bp_babord,                            --    conduit_end.bp_babord
			BP_Tribord => avalon_bouton_0_conduit_end_bp_tribord,                           --               .bp_tribord
			BP_STBY    => avalon_bouton_0_conduit_end_bp_stby,                              --               .bp_stby
			ledBabord  => avalon_bouton_0_conduit_end_ledbabord,                            --               .ledbabord
			ledTribord => avalon_bouton_0_conduit_end_ledtribord,                           --               .ledtribord
			ledSTBY    => avalon_bouton_0_conduit_end_ledstby,                              --               .ledstby
			out_bip    => avalon_bouton_0_conduit_end_out_bip                               --               .out_bip
		);

	avalon_verin_0 : component avalon_verin
		port map (
			write_data_i => mm_interconnect_0_avalon_verin_0_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			read_data_o  => mm_interconnect_0_avalon_verin_0_avalon_slave_0_readdata,  --               .readdata
			address_i    => mm_interconnect_0_avalon_verin_0_avalon_slave_0_address,   --               .address
			write_i      => mm_interconnect_0_avalon_verin_0_avalon_slave_0_write,     --               .write
			read_i       => mm_interconnect_0_avalon_verin_0_avalon_slave_0_read,      --               .read
			sck_o        => avalon_verin_0_conduit_end_sck_o,                          --    conduit_end.sck_o
			pwm_o        => avalon_verin_0_conduit_end_pwm_o,                          --               .pwm_o
			sens_o       => avalon_verin_0_conduit_end_sens_o,                         --               .sens_o
			miso_i       => avalon_verin_0_conduit_end_miso_i,                         --               .miso_i
			cs_n_o       => avalon_verin_0_conduit_end_cs_n_o,                         --               .cs_n_o
			clk_i        => clk_clk,                                                   --     clock_sink.clk
			arst_i       => rst_controller_reset_out_reset                             --     reset_sink.reset
		);

	boutons : component mon_sopc_boutons
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_boutons_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_boutons_s1_readdata,    --                    .readdata
			in_port  => boutons_external_connection_export        -- external_connection.export
		);

	jtag_uart_0 : component mon_sopc_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	leds : component mon_sopc_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	nios2_gen2_0 : component mon_sopc_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	ram : component mon_sopc_ram
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	test_anemo_0 : component avalon_gestion_anemometre
		port map (
			chipselect         => mm_interconnect_0_test_anemo_0_avalon_slave_0_chipselect,      -- avalon_slave_0.chipselect
			write_n            => mm_interconnect_0_test_anemo_0_avalon_slave_0_write_ports_inv, --               .write_n
			writedata          => mm_interconnect_0_test_anemo_0_avalon_slave_0_writedata,       --               .writedata
			readdata           => mm_interconnect_0_test_anemo_0_avalon_slave_0_readdata,        --               .readdata
			address            => mm_interconnect_0_test_anemo_0_avalon_slave_0_address,         --               .address
			reset_n            => rst_controller_reset_out_reset_ports_inv,                      --          reset.reset_n
			clk_50M            => clk_clk,                                                       --     clock_sink.clk
			in_freq_anemometre => test_anemo_0_conduit_end_beginbursttransfer                    --    conduit_end.beginbursttransfer
		);

	test_pwm_0 : component avalon_pwm
		port map (
			clk        => clk_clk,                                                     --          clock.clk
			chipselect => mm_interconnect_0_test_pwm_0_avalon_slave_0_chipselect,      -- avalon_slave_0.chipselect
			write_n    => mm_interconnect_0_test_pwm_0_avalon_slave_0_write_ports_inv, --               .write_n
			writedata  => mm_interconnect_0_test_pwm_0_avalon_slave_0_writedata,       --               .writedata
			readdata   => mm_interconnect_0_test_pwm_0_avalon_slave_0_readdata,        --               .readdata
			address    => mm_interconnect_0_test_pwm_0_avalon_slave_0_address,         --               .address
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --          reset.reset_n
			out_pwm    => test_pwm_0_conduit_end_writeresponsevalid_n                  --    conduit_end.writeresponsevalid_n
		);

	mm_interconnect_0 : component mon_sopc_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                     --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                            --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                        --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                         --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                               --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                           --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                              --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                          --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                        --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                     --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                 --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                        --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                    --                                         .readdata
			avalon_bouton_0_avalon_slave_0_address         => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_address,    --           avalon_bouton_0_avalon_slave_0.address
			avalon_bouton_0_avalon_slave_0_write           => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write,      --                                         .write
			avalon_bouton_0_avalon_slave_0_readdata        => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_readdata,   --                                         .readdata
			avalon_bouton_0_avalon_slave_0_writedata       => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_writedata,  --                                         .writedata
			avalon_bouton_0_avalon_slave_0_chipselect      => mm_interconnect_0_avalon_bouton_0_avalon_slave_0_chipselect, --                                         .chipselect
			avalon_verin_0_avalon_slave_0_address          => mm_interconnect_0_avalon_verin_0_avalon_slave_0_address,     --            avalon_verin_0_avalon_slave_0.address
			avalon_verin_0_avalon_slave_0_write            => mm_interconnect_0_avalon_verin_0_avalon_slave_0_write,       --                                         .write
			avalon_verin_0_avalon_slave_0_read             => mm_interconnect_0_avalon_verin_0_avalon_slave_0_read,        --                                         .read
			avalon_verin_0_avalon_slave_0_readdata         => mm_interconnect_0_avalon_verin_0_avalon_slave_0_readdata,    --                                         .readdata
			avalon_verin_0_avalon_slave_0_writedata        => mm_interconnect_0_avalon_verin_0_avalon_slave_0_writedata,   --                                         .writedata
			boutons_s1_address                             => mm_interconnect_0_boutons_s1_address,                        --                               boutons_s1.address
			boutons_s1_readdata                            => mm_interconnect_0_boutons_s1_readdata,                       --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			leds_s1_address                                => mm_interconnect_0_leds_s1_address,                           --                                  leds_s1.address
			leds_s1_write                                  => mm_interconnect_0_leds_s1_write,                             --                                         .write
			leds_s1_readdata                               => mm_interconnect_0_leds_s1_readdata,                          --                                         .readdata
			leds_s1_writedata                              => mm_interconnect_0_leds_s1_writedata,                         --                                         .writedata
			leds_s1_chipselect                             => mm_interconnect_0_leds_s1_chipselect,                        --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                         .debugaccess
			ram_s1_address                                 => mm_interconnect_0_ram_s1_address,                            --                                   ram_s1.address
			ram_s1_write                                   => mm_interconnect_0_ram_s1_write,                              --                                         .write
			ram_s1_readdata                                => mm_interconnect_0_ram_s1_readdata,                           --                                         .readdata
			ram_s1_writedata                               => mm_interconnect_0_ram_s1_writedata,                          --                                         .writedata
			ram_s1_byteenable                              => mm_interconnect_0_ram_s1_byteenable,                         --                                         .byteenable
			ram_s1_chipselect                              => mm_interconnect_0_ram_s1_chipselect,                         --                                         .chipselect
			ram_s1_clken                                   => mm_interconnect_0_ram_s1_clken,                              --                                         .clken
			test_anemo_0_avalon_slave_0_address            => mm_interconnect_0_test_anemo_0_avalon_slave_0_address,       --              test_anemo_0_avalon_slave_0.address
			test_anemo_0_avalon_slave_0_write              => mm_interconnect_0_test_anemo_0_avalon_slave_0_write,         --                                         .write
			test_anemo_0_avalon_slave_0_readdata           => mm_interconnect_0_test_anemo_0_avalon_slave_0_readdata,      --                                         .readdata
			test_anemo_0_avalon_slave_0_writedata          => mm_interconnect_0_test_anemo_0_avalon_slave_0_writedata,     --                                         .writedata
			test_anemo_0_avalon_slave_0_chipselect         => mm_interconnect_0_test_anemo_0_avalon_slave_0_chipselect,    --                                         .chipselect
			test_pwm_0_avalon_slave_0_address              => mm_interconnect_0_test_pwm_0_avalon_slave_0_address,         --                test_pwm_0_avalon_slave_0.address
			test_pwm_0_avalon_slave_0_write                => mm_interconnect_0_test_pwm_0_avalon_slave_0_write,           --                                         .write
			test_pwm_0_avalon_slave_0_readdata             => mm_interconnect_0_test_pwm_0_avalon_slave_0_readdata,        --                                         .readdata
			test_pwm_0_avalon_slave_0_writedata            => mm_interconnect_0_test_pwm_0_avalon_slave_0_writedata,       --                                         .writedata
			test_pwm_0_avalon_slave_0_chipselect           => mm_interconnect_0_test_pwm_0_avalon_slave_0_chipselect       --                                         .chipselect
		);

	irq_mapper : component mon_sopc_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_test_pwm_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_test_pwm_0_avalon_slave_0_write;

	mm_interconnect_0_test_anemo_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_test_anemo_0_avalon_slave_0_write;

	mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_avalon_bouton_0_avalon_slave_0_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of mon_sopc
