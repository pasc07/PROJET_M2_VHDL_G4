-- sopc_be.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sopc_be_1 is
	port (
		avalon_pwm_0_conduit_end_response   : out std_logic;                                       --     avalon_pwm_0_conduit_end.response
		clk_clk                             : in  std_logic                    := '0';             --                          clk.clk
		gpio_in_external_connection_export  : in  std_logic_vector(7 downto 0) := (others => '0'); --  gpio_in_external_connection.export
		gpio_out_external_connection_export : out std_logic_vector(7 downto 0);                    -- gpio_out_external_connection.export
		uart_external_connection_rxd        : in  std_logic                    := '0';             --     uart_external_connection.rxd
		uart_external_connection_txd        : out std_logic                                        --                             .txd
	);
end entity sopc_be_1;

architecture rtl of sopc_be_1 is
	component avalon_pwm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			out_pwm    : out std_logic                                         -- response
		);
	end component avalon_pwm;

	component sopc_be_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component sopc_be_cpu;

	component sopc_be_gpio_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component sopc_be_gpio_in;

	component sopc_be_gpio_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component sopc_be_gpio_out;

	component sopc_be_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sopc_be_jtag;

	component sopc_be_onchip_memory is
		port (
			clk        : in  std_logic                       := 'X';             -- clk
			address    : in  std_logic_vector(8 downto 0)    := (others => 'X'); -- address
			clken      : in  std_logic                       := 'X';             -- clken
			chipselect : in  std_logic                       := 'X';             -- chipselect
			write      : in  std_logic                       := 'X';             -- write
			readdata   : out std_logic_vector(1023 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(1023 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(127 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                       := 'X';             -- reset
			reset_req  : in  std_logic                       := 'X';             -- reset_req
			freeze     : in  std_logic                       := 'X'              -- freeze
		);
	end component sopc_be_onchip_memory;

	component sopc_be_sysid_1 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component sopc_be_sysid_1;

	component sopc_be_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component sopc_be_uart;

	component sopc_be_mm_interconnect_0 is
		port (
			clk_clk_clk                            : in  std_logic                       := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset  : in  std_logic                       := 'X';             -- reset
			jtag_reset_reset_bridge_in_reset_reset : in  std_logic                       := 'X';             -- reset
			cpu_data_master_address                : in  std_logic_vector(17 downto 0)   := (others => 'X'); -- address
			cpu_data_master_waitrequest            : out std_logic;                                          -- waitrequest
			cpu_data_master_byteenable             : in  std_logic_vector(3 downto 0)    := (others => 'X'); -- byteenable
			cpu_data_master_read                   : in  std_logic                       := 'X';             -- read
			cpu_data_master_readdata               : out std_logic_vector(31 downto 0);                      -- readdata
			cpu_data_master_write                  : in  std_logic                       := 'X';             -- write
			cpu_data_master_writedata              : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- writedata
			cpu_data_master_debugaccess            : in  std_logic                       := 'X';             -- debugaccess
			cpu_instruction_master_address         : in  std_logic_vector(17 downto 0)   := (others => 'X'); -- address
			cpu_instruction_master_waitrequest     : out std_logic;                                          -- waitrequest
			cpu_instruction_master_read            : in  std_logic                       := 'X';             -- read
			cpu_instruction_master_readdata        : out std_logic_vector(31 downto 0);                      -- readdata
			avalon_pwm_0_avalon_slave_0_address    : out std_logic_vector(1 downto 0);                       -- address
			avalon_pwm_0_avalon_slave_0_write      : out std_logic;                                          -- write
			avalon_pwm_0_avalon_slave_0_readdata   : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			avalon_pwm_0_avalon_slave_0_writedata  : out std_logic_vector(31 downto 0);                      -- writedata
			avalon_pwm_0_avalon_slave_0_chipselect : out std_logic;                                          -- chipselect
			cpu_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                       -- address
			cpu_debug_mem_slave_write              : out std_logic;                                          -- write
			cpu_debug_mem_slave_read               : out std_logic;                                          -- read
			cpu_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                      -- writedata
			cpu_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                       -- byteenable
			cpu_debug_mem_slave_waitrequest        : in  std_logic                       := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess        : out std_logic;                                          -- debugaccess
			gpio_in_s1_address                     : out std_logic_vector(1 downto 0);                       -- address
			gpio_in_s1_readdata                    : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			gpio_out_s1_address                    : out std_logic_vector(1 downto 0);                       -- address
			gpio_out_s1_write                      : out std_logic;                                          -- write
			gpio_out_s1_readdata                   : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			gpio_out_s1_writedata                  : out std_logic_vector(31 downto 0);                      -- writedata
			gpio_out_s1_chipselect                 : out std_logic;                                          -- chipselect
			jtag_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                       -- address
			jtag_avalon_jtag_slave_write           : out std_logic;                                          -- write
			jtag_avalon_jtag_slave_read            : out std_logic;                                          -- read
			jtag_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                      -- writedata
			jtag_avalon_jtag_slave_waitrequest     : in  std_logic                       := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect      : out std_logic;                                          -- chipselect
			onchip_memory_s1_address               : out std_logic_vector(8 downto 0);                       -- address
			onchip_memory_s1_write                 : out std_logic;                                          -- write
			onchip_memory_s1_readdata              : in  std_logic_vector(1023 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata             : out std_logic_vector(1023 downto 0);                    -- writedata
			onchip_memory_s1_byteenable            : out std_logic_vector(127 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect            : out std_logic;                                          -- chipselect
			onchip_memory_s1_clken                 : out std_logic;                                          -- clken
			sysid_1_control_slave_address          : out std_logic_vector(0 downto 0);                       -- address
			sysid_1_control_slave_readdata         : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- readdata
			uart_s1_address                        : out std_logic_vector(2 downto 0);                       -- address
			uart_s1_write                          : out std_logic;                                          -- write
			uart_s1_read                           : out std_logic;                                          -- read
			uart_s1_readdata                       : in  std_logic_vector(15 downto 0)   := (others => 'X'); -- readdata
			uart_s1_writedata                      : out std_logic_vector(15 downto 0);                      -- writedata
			uart_s1_begintransfer                  : out std_logic;                                          -- begintransfer
			uart_s1_chipselect                     : out std_logic                                           -- chipselect
		);
	end component sopc_be_mm_interconnect_0;

	component sopc_be_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sopc_be_irq_mapper;

	component sopc_be_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sopc_be_rst_controller;

	component sopc_be_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sopc_be_rst_controller_001;

	signal cpu_debug_reset_request_reset                                 : std_logic;                       -- cpu:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0);   -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                       -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                       -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(17 downto 0);   -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);    -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                       -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                         : std_logic;                       -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0);   -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0);   -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                       -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(17 downto 0);   -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                       -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect           : std_logic;                       -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0);   -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest          : std_logic;                       -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);    -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read                 : std_logic;                       -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write                : std_logic;                       -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0);   -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_chipselect      : std_logic;                       -- mm_interconnect_0:avalon_pwm_0_avalon_slave_0_chipselect -> avalon_pwm_0:chipselect
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_readdata        : std_logic_vector(31 downto 0);   -- avalon_pwm_0:readdata -> mm_interconnect_0:avalon_pwm_0_avalon_slave_0_readdata
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_address         : std_logic_vector(1 downto 0);    -- mm_interconnect_0:avalon_pwm_0_avalon_slave_0_address -> avalon_pwm_0:address
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write           : std_logic;                       -- mm_interconnect_0:avalon_pwm_0_avalon_slave_0_write -> mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write:in
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_writedata       : std_logic_vector(31 downto 0);   -- mm_interconnect_0:avalon_pwm_0_avalon_slave_0_writedata -> avalon_pwm_0:writedata
	signal mm_interconnect_0_sysid_1_control_slave_readdata              : std_logic_vector(31 downto 0);   -- sysid_1:readdata -> mm_interconnect_0:sysid_1_control_slave_readdata
	signal mm_interconnect_0_sysid_1_control_slave_address               : std_logic_vector(0 downto 0);    -- mm_interconnect_0:sysid_1_control_slave_address -> sysid_1:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0);   -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                       -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                       -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);    -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                       -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);    -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                       -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0);   -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                 : std_logic;                       -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                   : std_logic_vector(1023 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                    : std_logic_vector(8 downto 0);    -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                 : std_logic_vector(127 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                      : std_logic;                       -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                  : std_logic_vector(1023 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                      : std_logic;                       -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_uart_s1_chipselect                          : std_logic;                       -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                            : std_logic_vector(15 downto 0);   -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                             : std_logic_vector(2 downto 0);    -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                                : std_logic;                       -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer                       : std_logic;                       -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                               : std_logic;                       -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                           : std_logic_vector(15 downto 0);   -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal mm_interconnect_0_gpio_out_s1_chipselect                      : std_logic;                       -- mm_interconnect_0:gpio_out_s1_chipselect -> gpio_out:chipselect
	signal mm_interconnect_0_gpio_out_s1_readdata                        : std_logic_vector(31 downto 0);   -- gpio_out:readdata -> mm_interconnect_0:gpio_out_s1_readdata
	signal mm_interconnect_0_gpio_out_s1_address                         : std_logic_vector(1 downto 0);    -- mm_interconnect_0:gpio_out_s1_address -> gpio_out:address
	signal mm_interconnect_0_gpio_out_s1_write                           : std_logic;                       -- mm_interconnect_0:gpio_out_s1_write -> mm_interconnect_0_gpio_out_s1_write:in
	signal mm_interconnect_0_gpio_out_s1_writedata                       : std_logic_vector(31 downto 0);   -- mm_interconnect_0:gpio_out_s1_writedata -> gpio_out:writedata
	signal mm_interconnect_0_gpio_in_s1_readdata                         : std_logic_vector(31 downto 0);   -- gpio_in:readdata -> mm_interconnect_0:gpio_in_s1_readdata
	signal mm_interconnect_0_gpio_in_s1_address                          : std_logic_vector(1 downto 0);    -- mm_interconnect_0:gpio_in_s1_address -> gpio_in:address
	signal irq_mapper_receiver0_irq                                      : std_logic;                       -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                       -- uart:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0);   -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                : std_logic;                       -- rst_controller:reset_out -> [mm_interconnect_0:jtag_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                       -- rst_controller:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                       -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                       -- rst_controller_001:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv       : std_logic;                       -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv      : std_logic;                       -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write_ports_inv : std_logic;                       -- mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write:inv -> avalon_pwm_0:write_n
	signal mm_interconnect_0_uart_s1_read_ports_inv                      : std_logic;                       -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv                     : std_logic;                       -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal mm_interconnect_0_gpio_out_s1_write_ports_inv                 : std_logic;                       -- mm_interconnect_0_gpio_out_s1_write:inv -> gpio_out:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                       -- rst_controller_reset_out_reset:inv -> [avalon_pwm_0:reset_n, gpio_in:reset_n, gpio_out:reset_n, jtag:rst_n, sysid_1:reset_n, uart:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                       -- rst_controller_001_reset_out_reset:inv -> cpu:reset_n

begin

	avalon_pwm_0 : component avalon_pwm
		port map (
			clk        => clk_clk,                                                       --          clock.clk
			chipselect => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_chipselect,      -- avalon_slave_0.chipselect
			write_n    => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write_ports_inv, --               .write_n
			writedata  => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_writedata,       --               .writedata
			readdata   => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_readdata,        --               .readdata
			address    => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_address,         --               .address
			reset_n    => rst_controller_reset_out_reset_ports_inv,                      --          reset.reset_n
			out_pwm    => avalon_pwm_0_conduit_end_response                              --    conduit_end.response
		);

	cpu : component sopc_be_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	gpio_in : component sopc_be_gpio_in
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_gpio_in_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_gpio_in_s1_readdata,    --                    .readdata
			in_port  => gpio_in_external_connection_export        -- external_connection.export
		);

	gpio_out : component sopc_be_gpio_out
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_gpio_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_gpio_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_gpio_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_gpio_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_gpio_out_s1_readdata,        --                    .readdata
			out_port   => gpio_out_external_connection_export            -- external_connection.export
		);

	jtag : component sopc_be_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	onchip_memory : component sopc_be_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	sysid_1 : component sopc_be_sysid_1
		port map (
			clock    => clk_clk,                                            --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --         reset.reset_n
			readdata => mm_interconnect_0_sysid_1_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_1_control_slave_address(0)  --              .address
		);

	uart : component sopc_be_uart
		port map (
			clk           => clk_clk,                                   --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => uart_external_connection_rxd,              -- external_connection.export
			txd           => uart_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver1_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component sopc_be_mm_interconnect_0
		port map (
			clk_clk_clk                            => clk_clk,                                                  --                          clk_clk.clk
			cpu_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                       --  cpu_reset_reset_bridge_in_reset.reset
			jtag_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                           -- jtag_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                => cpu_data_master_address,                                  --                  cpu_data_master.address
			cpu_data_master_waitrequest            => cpu_data_master_waitrequest,                              --                                 .waitrequest
			cpu_data_master_byteenable             => cpu_data_master_byteenable,                               --                                 .byteenable
			cpu_data_master_read                   => cpu_data_master_read,                                     --                                 .read
			cpu_data_master_readdata               => cpu_data_master_readdata,                                 --                                 .readdata
			cpu_data_master_write                  => cpu_data_master_write,                                    --                                 .write
			cpu_data_master_writedata              => cpu_data_master_writedata,                                --                                 .writedata
			cpu_data_master_debugaccess            => cpu_data_master_debugaccess,                              --                                 .debugaccess
			cpu_instruction_master_address         => cpu_instruction_master_address,                           --           cpu_instruction_master.address
			cpu_instruction_master_waitrequest     => cpu_instruction_master_waitrequest,                       --                                 .waitrequest
			cpu_instruction_master_read            => cpu_instruction_master_read,                              --                                 .read
			cpu_instruction_master_readdata        => cpu_instruction_master_readdata,                          --                                 .readdata
			avalon_pwm_0_avalon_slave_0_address    => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_address,    --      avalon_pwm_0_avalon_slave_0.address
			avalon_pwm_0_avalon_slave_0_write      => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write,      --                                 .write
			avalon_pwm_0_avalon_slave_0_readdata   => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_readdata,   --                                 .readdata
			avalon_pwm_0_avalon_slave_0_writedata  => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_writedata,  --                                 .writedata
			avalon_pwm_0_avalon_slave_0_chipselect => mm_interconnect_0_avalon_pwm_0_avalon_slave_0_chipselect, --                                 .chipselect
			cpu_debug_mem_slave_address            => mm_interconnect_0_cpu_debug_mem_slave_address,            --              cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write              => mm_interconnect_0_cpu_debug_mem_slave_write,              --                                 .write
			cpu_debug_mem_slave_read               => mm_interconnect_0_cpu_debug_mem_slave_read,               --                                 .read
			cpu_debug_mem_slave_readdata           => mm_interconnect_0_cpu_debug_mem_slave_readdata,           --                                 .readdata
			cpu_debug_mem_slave_writedata          => mm_interconnect_0_cpu_debug_mem_slave_writedata,          --                                 .writedata
			cpu_debug_mem_slave_byteenable         => mm_interconnect_0_cpu_debug_mem_slave_byteenable,         --                                 .byteenable
			cpu_debug_mem_slave_waitrequest        => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,        --                                 .waitrequest
			cpu_debug_mem_slave_debugaccess        => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,        --                                 .debugaccess
			gpio_in_s1_address                     => mm_interconnect_0_gpio_in_s1_address,                     --                       gpio_in_s1.address
			gpio_in_s1_readdata                    => mm_interconnect_0_gpio_in_s1_readdata,                    --                                 .readdata
			gpio_out_s1_address                    => mm_interconnect_0_gpio_out_s1_address,                    --                      gpio_out_s1.address
			gpio_out_s1_write                      => mm_interconnect_0_gpio_out_s1_write,                      --                                 .write
			gpio_out_s1_readdata                   => mm_interconnect_0_gpio_out_s1_readdata,                   --                                 .readdata
			gpio_out_s1_writedata                  => mm_interconnect_0_gpio_out_s1_writedata,                  --                                 .writedata
			gpio_out_s1_chipselect                 => mm_interconnect_0_gpio_out_s1_chipselect,                 --                                 .chipselect
			jtag_avalon_jtag_slave_address         => mm_interconnect_0_jtag_avalon_jtag_slave_address,         --           jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write           => mm_interconnect_0_jtag_avalon_jtag_slave_write,           --                                 .write
			jtag_avalon_jtag_slave_read            => mm_interconnect_0_jtag_avalon_jtag_slave_read,            --                                 .read
			jtag_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                                 .readdata
			jtag_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                                 .writedata
			jtag_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                                 .waitrequest
			jtag_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      --                                 .chipselect
			onchip_memory_s1_address               => mm_interconnect_0_onchip_memory_s1_address,               --                 onchip_memory_s1.address
			onchip_memory_s1_write                 => mm_interconnect_0_onchip_memory_s1_write,                 --                                 .write
			onchip_memory_s1_readdata              => mm_interconnect_0_onchip_memory_s1_readdata,              --                                 .readdata
			onchip_memory_s1_writedata             => mm_interconnect_0_onchip_memory_s1_writedata,             --                                 .writedata
			onchip_memory_s1_byteenable            => mm_interconnect_0_onchip_memory_s1_byteenable,            --                                 .byteenable
			onchip_memory_s1_chipselect            => mm_interconnect_0_onchip_memory_s1_chipselect,            --                                 .chipselect
			onchip_memory_s1_clken                 => mm_interconnect_0_onchip_memory_s1_clken,                 --                                 .clken
			sysid_1_control_slave_address          => mm_interconnect_0_sysid_1_control_slave_address,          --            sysid_1_control_slave.address
			sysid_1_control_slave_readdata         => mm_interconnect_0_sysid_1_control_slave_readdata,         --                                 .readdata
			uart_s1_address                        => mm_interconnect_0_uart_s1_address,                        --                          uart_s1.address
			uart_s1_write                          => mm_interconnect_0_uart_s1_write,                          --                                 .write
			uart_s1_read                           => mm_interconnect_0_uart_s1_read,                           --                                 .read
			uart_s1_readdata                       => mm_interconnect_0_uart_s1_readdata,                       --                                 .readdata
			uart_s1_writedata                      => mm_interconnect_0_uart_s1_writedata,                      --                                 .writedata
			uart_s1_begintransfer                  => mm_interconnect_0_uart_s1_begintransfer,                  --                                 .begintransfer
			uart_s1_chipselect                     => mm_interconnect_0_uart_s1_chipselect                      --                                 .chipselect
		);

	irq_mapper : component sopc_be_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component sopc_be_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,      -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component sopc_be_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,          -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_avalon_pwm_0_avalon_slave_0_write;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	mm_interconnect_0_gpio_out_s1_write_ports_inv <= not mm_interconnect_0_gpio_out_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of sopc_be
